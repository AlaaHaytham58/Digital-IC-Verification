`ifndef ALU_env_SVH
`define ALU_env_SVH
`include "uvm_macros.svh"

`include  "alu_agent.svh"

import uvm_pkg::*;
class alu_env extends uvm_env;
    alu_agent agent;
    `uvm_component_utils(alu_env)
    function new(string name="alu_env",uvm_component parent =null);
        super.new(name,parent);
    endfunction
    function void buildphase(uvm_phase phase);
     super.build_phase(phase);
     `uvm_info("KAMONNNNA","alu env build phase",UVM_LOW)
    endfunction
endclass
`endif
package alu_pkg;
`include "alu_transaction.svh"
`include "alu_test.svh"
endpackage
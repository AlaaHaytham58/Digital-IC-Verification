interface alu_if;
 logic clk;
 logic rst;
 logic [3:0]a;
 logic[3:0]b;
 logic [1:0]op;
 logic [3:0]result;
endinterface